/*

 */
`default_nettype none
`timescale 1ns/1ps
module test_sdd(
           input wire clk_25mhz,
           inout wire [GPIO_NR -1:0] gpio,
           output wire [24:21] gn,
           output wire [24:21] gp
       );

//localparam SYSTEM_CLK = 110_000_000;
localparam SYSTEM_CLK = 80_000_000;
localparam GPIO_NR = 8;
 /* gpio */
 reg  [GPIO_NR -1:0] gpio_output_en;
 wire [GPIO_NR -1:0] gpio_in;
 reg  [GPIO_NR -1:0] gpio_output_val;

wire [31:0] mem_din;

 wire gpio_output_wr;
 wire gpio_output_val_wr;
 wire gpio_output_en_wr;

 /* input */
 assign gpio_in = gpio;

 /* output */
 genvar i;
 generate
   for (i = 0; i < GPIO_NR; i = i +1) begin
     assign gpio[i] = gpio_output_en[i] ? gpio_output_val[i] : 1'bz;
   end
 endgenerate

 always @(posedge clk) begin
   if (!resetn) begin
     gpio_output_en  <=  0;  // default all is input pin
     gpio_output_val <=  0;  // digilent led 0: off 1:0
   end else begin
     gpio_output_val <= gpio_output_val_wr ? mem_din[GPIO_NR -1:0] : gpio_output_val;
     gpio_output_en  <= gpio_output_en_wr  ? mem_din[GPIO_NR -1:0] : gpio_output_en;
   end
 end

// reset
reg [15:0] reset_cnt = 0;
wire resetn = 0;
always @(posedge clk) begin
    if (reset_cnt == 0) begin
        resetn <= 1;
    end else begin
        resetn <= 0;
    end
    reset_cnt <= reset_cnt + {14'b0, !resetn};
end

//wire clk = clk_25mhz;
wire clk;
pll #(SYSTEM_CLK/1_000_000) pll_i(clk_25mhz, clk);

wire   oled_cs;
wire   oled_mosi;
wire   oled_sck;
wire   oled_dc;
wire   oled_rst;
wire   oled_vccen;
wire   oled_pmoden;
reg [7:0]    oled_x_dc;
reg [7:0]    oled_y_data;
reg [15:0]   oled_rgb;
reg          oled_strobe;
reg          oled_setpixel_raw8tx;

wire         oled_ready;
wire         oled_valid;
assign gn[24] = oled_cs;
assign gn[23] = oled_mosi;
assign gn[21] = oled_sck;

assign gp[24] = oled_dc;
assign gp[23] = oled_rst;
assign gp[22] = oled_vccen;
assign gp[21] = oled_pmoden;

sdd1331_gen_pattern ssd_clk(
           .clk(clk),
           .out_hcnt(oled_x_dc),
           .out_vcnt(oled_y_data),
           .rgb(oled_rgb),
           .rst(~resetn)
       );


oled_ssd1331 #(.SYSTEM_CLK(SYSTEM_CLK))
             oled_ssd1331_i(
                 .clk(clk),
                 .resetn(resetn),
                 .oled_rst(oled_rst),
                 .strobe(oled_strobe),
                 .setpixel_raw8tx(oled_setpixel_raw8tx),
                 .x_dc(oled_x_dc),
                 .y_data(oled_y_data),
                 .rgb(oled_rgb),
                 .ready(oled_ready),
                 .valid(oled_valid),
                 .spi_cs(oled_cs),
                 .spi_dc(oled_dc),
                 .spi_mosi(oled_mosi),
                 .spi_sck(oled_sck),
                 .vccen(oled_vccen),
                 .pmoden(oled_pmoden)
             );


endmodule

    /*
     * Do not edit this file, it was generated by gen_pll.sh
     *
     *   FPGA kind      : ECP5
     *   Input frequency: 25 MHz
     */

    module pll #(
        parameter freq = 40
    ) (
        input wire pclk,
        output wire clk
    );
(* ICP_CURRENT="12" *) (* LPF_RESISTOR="8" *) (* MFG_ENABLE_FILTEROPAMP="1" *) (* MFG_GMCREF_SEL="2" *)
EHXPLLL pll_i (
            .RST(1'b0),
            .STDBY(1'b0),
            .CLKI(pclk),
            .CLKOP(clk),
            .CLKFB(clk),
            .CLKINTFB(),
            .PHASESEL0(1'b0),
            .PHASESEL1(1'b0),
            .PHASEDIR(1'b1),
            .PHASESTEP(1'b1),
            .PHASELOADREG(1'b1),
            .PLLWAKESYNC(1'b0),
            .ENCLKOP(1'b0)
        );
defparam pll_i.PLLRST_ENA = "DISABLED";
defparam pll_i.INTFB_WAKE = "DISABLED";
defparam pll_i.STDBY_ENABLE = "DISABLED";
defparam pll_i.DPHASE_SOURCE = "DISABLED";
defparam pll_i.OUTDIVIDER_MUXA = "DIVA";
defparam pll_i.OUTDIVIDER_MUXB = "DIVB";
defparam pll_i.OUTDIVIDER_MUXC = "DIVC";
defparam pll_i.OUTDIVIDER_MUXD = "DIVD";
defparam pll_i.CLKOP_ENABLE = "ENABLED";
defparam pll_i.CLKOP_FPHASE = 0;
defparam pll_i.FEEDBK_PATH = "CLKOP";
generate
    case(freq)
        16: begin
            defparam pll_i.CLKI_DIV=8;
            defparam pll_i.CLKOP_DIV=38;
            defparam pll_i.CLKOP_CPHASE=18;
            defparam pll_i.CLKFB_DIV=5;
        end
        20: begin
            defparam pll_i.CLKI_DIV=5;
            defparam pll_i.CLKOP_DIV=30;
            defparam pll_i.CLKOP_CPHASE=15;
            defparam pll_i.CLKFB_DIV=4;
        end
        24: begin
            defparam pll_i.CLKI_DIV=1;
            defparam pll_i.CLKOP_DIV=24;
            defparam pll_i.CLKOP_CPHASE=11;
            defparam pll_i.CLKFB_DIV=1;
        end
        25: begin
            defparam pll_i.CLKI_DIV=1;
            defparam pll_i.CLKOP_DIV=24;
            defparam pll_i.CLKOP_CPHASE=11;
            defparam pll_i.CLKFB_DIV=1;
        end
        30: begin
            defparam pll_i.CLKI_DIV=5;
            defparam pll_i.CLKOP_DIV=20;
            defparam pll_i.CLKOP_CPHASE=9;
            defparam pll_i.CLKFB_DIV=6;
        end
        35: begin
            defparam pll_i.CLKI_DIV=5;
            defparam pll_i.CLKOP_DIV=17;
            defparam pll_i.CLKOP_CPHASE=8;
            defparam pll_i.CLKFB_DIV=7;
        end
        40: begin
            defparam pll_i.CLKI_DIV=5;
            defparam pll_i.CLKOP_DIV=15;
            defparam pll_i.CLKOP_CPHASE=7;
            defparam pll_i.CLKFB_DIV=8;
        end
        45: begin
            defparam pll_i.CLKI_DIV=5;
            defparam pll_i.CLKOP_DIV=13;
            defparam pll_i.CLKOP_CPHASE=6;
            defparam pll_i.CLKFB_DIV=9;
        end
        48: begin
            defparam pll_i.CLKI_DIV=8;
            defparam pll_i.CLKOP_DIV=13;
            defparam pll_i.CLKOP_CPHASE=6;
            defparam pll_i.CLKFB_DIV=15;
        end
        50: begin
            defparam pll_i.CLKI_DIV=1;
            defparam pll_i.CLKOP_DIV=12;
            defparam pll_i.CLKOP_CPHASE=5;
            defparam pll_i.CLKFB_DIV=2;
        end
        55: begin
            defparam pll_i.CLKI_DIV=5;
            defparam pll_i.CLKOP_DIV=11;
            defparam pll_i.CLKOP_CPHASE=5;
            defparam pll_i.CLKFB_DIV=11;
        end
        60: begin
            defparam pll_i.CLKI_DIV=5;
            defparam pll_i.CLKOP_DIV=10;
            defparam pll_i.CLKOP_CPHASE=4;
            defparam pll_i.CLKFB_DIV=12;
        end
        65: begin
            defparam pll_i.CLKI_DIV=5;
            defparam pll_i.CLKOP_DIV=9;
            defparam pll_i.CLKOP_CPHASE=4;
            defparam pll_i.CLKFB_DIV=13;
        end
        66: begin
            defparam pll_i.CLKI_DIV=8;
            defparam pll_i.CLKOP_DIV=9;
            defparam pll_i.CLKOP_CPHASE=4;
            defparam pll_i.CLKFB_DIV=21;
        end
        70: begin
            defparam pll_i.CLKI_DIV=5;
            defparam pll_i.CLKOP_DIV=9;
            defparam pll_i.CLKOP_CPHASE=4;
            defparam pll_i.CLKFB_DIV=14;
        end
        75: begin
            defparam pll_i.CLKI_DIV=1;
            defparam pll_i.CLKOP_DIV=8;
            defparam pll_i.CLKOP_CPHASE=4;
            defparam pll_i.CLKFB_DIV=3;
        end
        80: begin
            defparam pll_i.CLKI_DIV=5;
            defparam pll_i.CLKOP_DIV=7;
            defparam pll_i.CLKOP_CPHASE=3;
            defparam pll_i.CLKFB_DIV=16;
        end
        85: begin
            defparam pll_i.CLKI_DIV=5;
            defparam pll_i.CLKOP_DIV=7;
            defparam pll_i.CLKOP_CPHASE=3;
            defparam pll_i.CLKFB_DIV=17;
        end
        90: begin
            defparam pll_i.CLKI_DIV=5;
            defparam pll_i.CLKOP_DIV=7;
            defparam pll_i.CLKOP_CPHASE=3;
            defparam pll_i.CLKFB_DIV=18;
        end
        95: begin
            defparam pll_i.CLKI_DIV=5;
            defparam pll_i.CLKOP_DIV=6;
            defparam pll_i.CLKOP_CPHASE=3;
            defparam pll_i.CLKFB_DIV=19;
        end
        100: begin
            defparam pll_i.CLKI_DIV=1;
            defparam pll_i.CLKOP_DIV=6;
            defparam pll_i.CLKOP_CPHASE=2;
            defparam pll_i.CLKFB_DIV=4;
        end
        105: begin
            defparam pll_i.CLKI_DIV=5;
            defparam pll_i.CLKOP_DIV=6;
            defparam pll_i.CLKOP_CPHASE=2;
            defparam pll_i.CLKFB_DIV=21;
        end
        110: begin
            defparam pll_i.CLKI_DIV=5;
            defparam pll_i.CLKOP_DIV=5;
            defparam pll_i.CLKOP_CPHASE=2;
            defparam pll_i.CLKFB_DIV=22;
        end
        115: begin
            defparam pll_i.CLKI_DIV=5;
            defparam pll_i.CLKOP_DIV=5;
            defparam pll_i.CLKOP_CPHASE=2;
            defparam pll_i.CLKFB_DIV=23;
        end
        120: begin
            defparam pll_i.CLKI_DIV=5;
            defparam pll_i.CLKOP_DIV=5;
            defparam pll_i.CLKOP_CPHASE=2;
            defparam pll_i.CLKFB_DIV=24;
        end
        125: begin
            defparam pll_i.CLKI_DIV=1;
            defparam pll_i.CLKOP_DIV=5;
            defparam pll_i.CLKOP_CPHASE=2;
            defparam pll_i.CLKFB_DIV=5;
        end
        130: begin
            defparam pll_i.CLKI_DIV=5;
            defparam pll_i.CLKOP_DIV=5;
            defparam pll_i.CLKOP_CPHASE=2;
            defparam pll_i.CLKFB_DIV=26;
        end
        135: begin
            defparam pll_i.CLKI_DIV=5;
            defparam pll_i.CLKOP_DIV=4;
            defparam pll_i.CLKOP_CPHASE=2;
            defparam pll_i.CLKFB_DIV=27;
        end
        140: begin
            defparam pll_i.CLKI_DIV=5;
            defparam pll_i.CLKOP_DIV=4;
            defparam pll_i.CLKOP_CPHASE=1;
            defparam pll_i.CLKFB_DIV=28;
        end
        default: UNKNOWN_FREQUENCY unknown_frequency();
    endcase
endgenerate
endmodule
